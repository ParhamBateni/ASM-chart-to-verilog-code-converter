library verilog;
use verilog.vl_types.all;
entity module2 is
    port(
        S               : in     vl_logic_vector(31 downto 0);
        output2         : out    vl_logic_vector(31 downto 0)
    );
end module2;
