library verilog;
use verilog.vl_types.all;
entity module8 is
    port(
        R1              : in     vl_logic_vector(31 downto 0);
        output8         : out    vl_logic_vector(31 downto 0)
    );
end module8;
