library verilog;
use verilog.vl_types.all;
entity module5 is
    port(
        i               : in     vl_logic_vector(31 downto 0);
        e               : in     vl_logic_vector(31 downto 0);
        output5         : out    vl_logic_vector(31 downto 0)
    );
end module5;
